`timescale 1ps/1ns
 module lab9()




 endmodule